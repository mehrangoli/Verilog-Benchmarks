/*
Author: Mehran Goli
Version: 1.0
Date: 17-8-2019
*/
module add(in1,in2,cin,cout,out);
	
	input  in1,in2,cin; 
	output cout,out; 
	
////////////////////////////////////////////////////////////////////////////////////////////

	assign {cout,out} = in1+in2+cin ;
/////////////////////////////////////////////////////////////////////////////////////////////////	

endmodule
